module Swiches_To_LEDs(
	input i_Switch_1,
	input i_Switch_2,
	input i_Switch_3,
	input i_Switch_4,
	output o_LED_1,
	output o_LED_2,
	output o_LED_3,
	output o_LED_4);
	
	assign i_Switch_1 = i_Switch_1;
	assign i_Switch_2 = i_Switch_2;
	assign i_Switch_3 = i_Switch_3;
	assign i_Switch_4 = i_Switch_4;
	
endmodule // Swiches_To_LEDs
	
	